module top #(RAM1_DATA_WIDTH = 32, RAM2_DATA_WIDTH = 16, ADDR_WIDTH = 4, DEPTH = 32) (a, Output,clk);

    //Mac1 and sram inputs

    input wire [7:0] ip_attr;
    input wire clk, rst, we, i_write;
    input wire [31:0] ram_1_data_in;
    input wire [ADDR_WIDTH-1:0] in_addr;
    input wire [RAM1_DATA_WIDTH-1:0] ram1_data_in;
    input wire [RAM2_DATA_WIDTH-1:0] ram2_data_in;

    //Mac1 output
    reg [15:0] mac_acc;
    //Ram1 and Ram2 inputs
    reg ram1clk;
    reg ram2clk;
    //Ram1 and Ram2 outputs
    reg [RAM1_DATA_WIDTH-1:0 ram1reg;
    reg [RAM2_DATA_WIDTH-1:0] ram2reg;

    //Instantiate clkdiv to reduce clkfreq by 4 times for Ram1 and to half the clkfreq for RAM2_DATA_WIDTH
    //So total 2 clkdiv modules
    clkdiv #(.DIVISOR(4)) clkdivram1 (
        .clock_in(clk),
        .clock_out(ram1clk)
        );

    clkdiv #(.DIVISOR(2)) clkdivram2 (
        .clock_in(clk),
        .clock_out(ram2clk)
        );

    





























// input wire a[31:0];
//
// input wire clk;
// output reg[8:0] Output;
//
//
// reg[7:0] a,b;
// reg[7:0] na =8'b00000000;;      //next address/class
// reg c =1'b0;          //class flag
// reg [7:0] c1,c2,c3,c4;
// reg [15:0] t;
// reg count;
//
//
//
//     sram1  sram_node (
//     .i_clk(clk),
//     .i_addr(node_addr),
//     .i_write(i_write),
//     .i_data(i_data),
//     .o_data(coeff)
// );
//
//     sram2  sram_child (
//     .i_clk(clk),
//     .i_addr(inputAddr),
//     .i_write(i_write),
//     .i_da(i_data),
//     .o_da(child)
// );
//     mac1 mac_i(.a(a),.b(b),.c3(c3),.rst(rst), .acc(acc) clk(clk));
//
//
// assign i_write=0;
// assign i_data=1;
//
//
// //always@(a)
// //c=0;
// while (c==0) begin
//
//
// begin
//     count=0;
//     inputAddr=na[7:0];
//     c1=coeff[32:24];c2=coeff[23:16];c3=coeff[15:8];c4=coeff[7:0];
//     always @ (clk) begin
//       if (count==0) begin
//       rst=1;
//       a = c1; b=a[23:16];
//       rst=0;
//       count= count+1;
//       end
//       if (count==1) begin
//       a = c2; b=a[15:8];
//       count= count+1;
//       if (count==2) begin
//       a = c3; b=a[7:0];
//       t=acc;
//       count= 0;
//     end
//
//
//
//   if  (t < c4)
//     begin
//         assign na=child[17:9];  //child address including the chld or class bit, so total 11+1=12 bits
//     end
//   else
//     begin
//         assign na=child[8:0];
//     end
//
//
//     if na[8]==1
//     begin
//       assign c=1;
//       Output=child;
//      end
// end



endmodule // top
